package Deserializer(
  mkSeserialize,
  ISeserializer(..),
  State(..)) 
  where

import ClkDivider
import State

serialize :: State -> Bit 8 -> Bit 1
serialize ftdiState dataReg =
    case ftdiState of
        START    -> 1'b0
        (DATA n) -> dataReg[0]
        _        -> 1'b1
-- serialize START _ = 1'b0
-- serialize (DATA n) data = data[n]
-- serialize _ _ = 1'b1

interface (ISeserializer :: # -> # -> *) clkFreq baudRate = 
  putBit8    :: (Bit 8) -> Action {-# always_enabled, always_ready #-}
  bitLineOut ::  Bit 1            {-# always_ready #-}

mkSeserialize :: Handle -> Module (IDeserializer clkFreq baudRate)
mkSeserialize fileHandle = do

  ftdiTxOut :: Wire(Bit 1) <- mkBypassWire
  dataReg  :: Reg(Bit 8) <- mkReg(0)
  ftdiState <- mkReg(IDLE)
  clkDivider :: (ClkDivider (TDiv clkFreq baudRate)) <- mkClkDivider fileHandle

  addRules $
    rules
      {-# ASSERT fire when enabled #-}
      "ADVANCE UART STATE WHEN NOT IDLE" : when 
        (ftdiState /= IDLE), 
        (clkDivider.isAdvancing) ==>
        do
          ftdiState := ftdiState' ftdiState

      {-# ASSERT fire when enabled #-}
      "BIT LINE" : when True ==>
        do
          ftdiTxOut := serialize ftdiState dataReg

  return $
    interface ISeserializer
    {putBit8  bit8Val = 
        clkDivider.reset
        dataReg := bit8Val 
        ftdiState := ftdiState' ftdiState
        when (ftdiState == IDLE)
    ;bitLineOut = ftdiTxOut
    }