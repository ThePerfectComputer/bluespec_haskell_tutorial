package Util(simulate_for) where

simulate_for :: (Bits a n, Arith a, Eq a) => Reg a -> Reg a -> Rules
simulate_for curr_cycle end_cycle =
  rules
    "count_cycle_rule": when True ==> action
      curr_cycle := curr_cycle + 1
      if curr_cycle == end_cycle
        then 
          $finish
        else
          $display "cycle = " curr_cycle
