-- TOPMODULE=mkTop make b_compile
package Top(mkClkDivider, ClkDivider(..)) where

data State = IDLE | START | DATA (UInt (TLog 8)) | PARITY | STOP
  deriving (Bits, Eq, FShow)

type FCLK = 25_000_000
type BAUD = 9_600

interface (ClkDivider :: # -> *) hi =
  {
  reset :: Action
  ;isAdvancing :: Bool
  ;isHalfCycle :: Bool
  }

mkClkDivider :: Handle -> Module (ClkDivider hi)
mkClkDivider fileHandle = do
    counter <- mkReg(0 :: UInt (TLog hi))   
    let hi_value :: UInt (TLog hi) = (fromInteger $ valueOf hi)
    let half_hi_value :: UInt (TLog hi) = (fromInteger $ valueOf (TDiv hi 2))

    let val :: Real = (fromInteger $ valueOf hi)
    let msg = "Clock Div Period : " + (realToString val)
    -- messageM msg

    hPutStr fileHandle msg
    hPutStr fileHandle genModuleName
    -- hClose fileHandle

    addRules $
      rules
        {-# ASSERT fire when enabled #-}
        {-# ASSERT no implicit conditions #-}
        "tick" : when True ==> action
          $display (counter)
          counter := if (counter == hi_value)
                    then 0
                    else counter + 1
    
    return $
      interface ClkDivider
        reset :: Action
        reset = do
          counter := 0

        isAdvancing :: Bool
        isAdvancing = (counter == hi_value)
        isHalfCycle = (counter == half_hi_value)

interface (IDeserializer :: # -> # -> *) clkFreq baudRate = 
  get         ::  Bit 8            {-# always_ready #-}
  putBitIn    :: (Bit 1) -> Action {-# always_enabled, always_ready #-}

mkDeserialize :: Handle -> Module (IDeserializer clkFreq baudRate)
mkDeserialize fileHandle = do
  -- figure out why changing to wire below doesn't work
  ftdiRxIn :: Wire(Bit 1) <- mkBypassWire
  shiftReg :: Reg(Bit 8) <- mkReg(0)
  ftdiState <- mkReg(IDLE)

  clkDivider :: (ClkDivider (TDiv clkFreq baudRate)) <- mkClkDivider fileHandle

  addRules $
    rules

      {-# ASSERT fire when enabled #-}
      when (ftdiState == IDLE), (ftdiRxIn == 0) ==>
        do
          clkDivider.reset
          ftdiState := START 

      {-# ASSERT fire when enabled #-}
      when (ftdiState == START), (clkDivider.isAdvancing) ==>
        do
          ftdiState := DATA(0)

      {-# ASSERT fire when enabled #-}
        when 
          DATA(n) <- ftdiState,
          n >= 0,
          n <= 7, 
          let sampleTrigger = clkDivider.isHalfCycle
            in sampleTrigger
          ==>
            do
              ftdiState := 
                if n == 7
                  then PARITY
                  else DATA(n + 1)
              shiftReg := ftdiRxIn ++ shiftReg[7:1]

      {-# ASSERT fire when enabled #-}
      when (ftdiState == PARITY), (clkDivider.isAdvancing) ==>
        do
          ftdiState := STOP

      {-# ASSERT fire when enabled #-}
      when (ftdiState == STOP), (clkDivider.isAdvancing) ==>
        do
          ftdiState := IDLE

  return $
    interface IDeserializer
    {get      = shiftReg when (ftdiState == STOP), (clkDivider.isAdvancing)
    ;putBitIn bit = ftdiRxIn := bit
    }

interface ITop = 
  ftdi_rxd    ::  Bit 1            {-# always_ready #-}
  led         ::  Bit 8            {-# always_ready #-}
  ftdi_txd    :: (Bit 1) -> Action {-# always_enabled, always_ready #-}

{-# properties mkTop={verilog} #-}
mkTop :: Module (ITop)
mkTop = do

  fileHandle <- openFile "compile.log" WriteMode 

  serializer :: (IDeserializer FCLK BAUD) <- mkDeserialize fileHandle
  ftdiBitIn  :: Wire(Bit 1)       <- mkBypassWire
  rxReg      :: Reg(Bit 8) <- mkReg(0)

  addRules $
    rules
      when True ==>
        rxReg := serializer.get
      
      when True ==>
        serializer.putBitIn ftdiBitIn

  return $
    interface ITop
    {ftdi_rxd = ftdiBitIn
    ;led = rxReg
    ;ftdi_txd bitIn = ftdiBitIn := bitIn}

mkSim :: Module Empty
mkSim = do
  -- count :: Reg(UInt 3) <- mkReg(0)
  count :: Reg(UInt 3) <- mkReg(0)
  addRules $
    rules
      "count" : when True ==> action
        count := unpack ((1'b1) ++ (pack count)[2:1])
        $display count
      "end sim" : when (count == 6) ==> action
        $finish

  return $
    interface Empty