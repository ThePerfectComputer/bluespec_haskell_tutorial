-- should spit out the following when compiled
-- Compilation message: "src/Top.bs", line 11, column 45:  valueOf (TLog TestVal) 4.0
package Top where

type TestVal = 9

mkTop :: Module Empty
mkTop =
  module
    let testVal :: Integer
        testVal  = valueOf (TLog TestVal)

    messageM $ " valueOf (TLog TestVal) " + (realToString $ fromInteger testVal)

    addRules $
      rules
        when True ==> action
          $finish
