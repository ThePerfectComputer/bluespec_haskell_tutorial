package Top where
import List
import GetPut

data RxState = Idle | Capturing | Done | Error 
                deriving(Bits, Eq, FShow)

interface (Counter :: # -> *) hi =
  reset :: Action
  isSaturated :: ActionValue Bool

mkCounter :: Module (Counter hi)
mkCounter = 
  module
    counter <- mkReg(0 :: UInt (TLog hi))   
    let hi_value :: UInt (TLog hi) = (fromInteger $ valueOf hi)

    rules
      "count" : when True ==> action
        $display (counter)
        counter := if (counter == hi_value) then 0 else (counter + 1)
        counter := case counter of
                     hi_value -> 0
                     _        -> counter + 1
    
    interface
      reset :: Action
      reset = do
        counter := 0
      isSaturated :: ActionValue Bool
      isSaturated = do
        return (counter == hi_value)

interface UartRx =
  put_rx_bit  :: (Bit 1) -> Action
  get_rx_char :: ActionValue Char

-- mkUartRx :: UInt 32 -> Module (UartRx)
-- mkUartRx interval = 
--   module
--     rx_in           :: Wire (Bit 1) <- mkWire
--     rx_in_previous  :: Reg  (Maybe (Bit 1)) <- mkReg (Invalid)
--     rx_captured     :: Wire (Maybe (Bit 1)) <- mkWire
--     thing <- mkReg(True)

--     -- let num = 3
--     -- let num_bits      =  log2 $ fromInteger interval
--     interval_counter  :: Reg(UInt 32)
--     interval_counter  <- mkReg(interval)

--     rx_state          :: Reg(RxState) <- mkReg(Idle)

--     rules
--       "register_rx" : when True ==> action
--         rx_in_previous  := Valid rx_in
--         rx_captured     := case (rx_in_previous, rx_in) of 
--                               (Valid 1, 1) -> Valid 1
--                               (Valid 0, 0) -> Valid 0
--                               (_,_)        -> Invalid

--       "value_captured":
--         when Valid 1 <- rx_captured
--           ==> action
--             thing := False

--     let get = do {return ('a' :: Char)}

--     interface 
--       get_rx_char :: ActionValue Char
--       get_rx_char = get

--       put_rx_bit :: (Bit 1) -> Action
--       put_rx_bit bit_val = do
--         rx_in := bit_val

mkTop :: Module (Empty)
mkTop = 
  module
    sync_regs <- replicateM 2 (mkReg (0 :: UInt 2))
    let list1 :: List (UInt 32)  = (map fromInteger (upto 1 4))
    let list2 :: List (UInt 32)  = (map fromInteger (upto 2 9))
    -- let list3 :: List (UInt 32, UInt 32) = zip list1 list2
    let list3 = zip list1 list2
    counter <- mkReg(0 :: UInt 32)

    rules
      "reg_chain" : when True ==> action
        (sync_regs !! 0) := readReg (sync_regs !! 1)
      "simulate" : when counter < 5 ==> action
        counter := counter + 1
        if counter == 1 then
          do
            $finish
        else action {}
        $display (fshow list3)
    -- return Empty

mkSim :: Module Empty
mkSim =
  module
    my_counter :: Counter(3) <- mkCounter
    cycle  <- mkReg(0 :: UInt 32)

    rules
      "incr cycle": when True ==> action
        cycle := cycle + 1
        $display "my_counter " my_counter.isSaturated

      "end sim": when (cycle == 6) ==> action
        $finish