package Top where

interface Blinky =
    led        :: Bit 8
  
{-# properties mkBlinky={alwaysReady} #-}
mkBlinky :: Module (Blinky)
mkBlinky = 
  module
    counter   <- mkReg(0 :: UInt 32)

    rules 
      "incr": when True ==> action
        counter := counter + 1

    interface
      led        = (pack counter)[29:22]

mkSim :: Module Empty
mkSim =
  module
    dut <- mkBlinky
    old_led_val <- mkReg(0 :: Bit 8)

    cycle  <- mkReg(0 :: UInt 32)
    alerts <- mkReg(0 :: UInt 32)

    rules
      "incr cycle": when True ==> action
        cycle := cycle + 1

      "follow led": when True ==> action
        old_led_val := dut.led

      "notify change": when (old_led_val /= dut.led) ==> action
        $display "cycle = " cycle
        $display "dut.led = " dut.led
        alerts := alerts + 1

      "end sim": when (alerts == 6) ==> action
        $finish