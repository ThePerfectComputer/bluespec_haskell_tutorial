-- Copyright (c) 2014-2020 Bluespec, Inc.  All Rights Reserved.

package Top where

mkTop :: Module Empty
mkTop =
  module
    addRules mkHelloRule

mkHelloRule :: Rules
mkHelloRule = 
    rules
      "rl_print_answer": when True ==> action
          $display "Hello World."
          $finish