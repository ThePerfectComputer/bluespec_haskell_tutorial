package Top where

mkTop :: Module Empty
mkTop = do
  return $ interface Empty { }
