package Top where

mkTop :: Module Empty
mkTop =
  module
    -- I'm not declaring types for the reg here, it can be inferred,
    -- and later we could have a language server that allows for inspection
    -- of inferred types
    -- cycle :: Reg(Int 16)
    cycle <- mkReg (negate 1)
    end_cycle <- mkReg 4

    addRules $ mkHelloRule <+> (simulate_for cycle end_cycle)
    -- addRules $ (simulate_for cycle end_cycle) <+> mkHelloRule

mkHelloRule :: Rules
mkHelloRule = 
    rules
      "rl_print_answer": when True ==> action
          $display "Hello World." $stime

simulate_for :: (Bits a n, Arith a, Eq a) => Reg a -> Reg a -> Rules
simulate_for curr_cycle end_cycle =
  rules
    "count_cycle_rule": when True ==> action
      curr_cycle := curr_cycle + 1
      if curr_cycle == end_cycle
        then 
          $finish
        else
          $display curr_cycle
