package Top where

import Util

data AluState = Add | Subtract | Multiply deriving(Bits, Eq, FShow)

mkTop :: Module Empty
mkTop =
  module
    -- allows us to run and end the simulation
    cycle <- mkReg 0
    end_cycle <- mkReg 4
    addRules (simulate_for cycle end_cycle)

    -- build what is basically an alu with a state register
    state :: Reg(AluState)
    state <- mkReg(Add)

    a :: Reg(Int 32)
    a <- mkReg 10

    b :: Reg(Int 32)
    b <- mkReg 12

    o :: Wire(Int 32)
    o <- mkWire

    rules
      "alu": when True ==> action
        o := 
          case state of
            Add      -> a + b
            Subtract -> a - b
            Multiply -> a * b

      "cycle_state": when True ==> action
        state :=
          case state of
            Add      -> Subtract
            Subtract -> Multiply
            Multiply -> Add
      
      "display": when True ==> action
        $display "alu.o = " o
        $display "state = " (fshow state)
      