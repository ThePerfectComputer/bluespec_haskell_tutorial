-- TOPMODULE=mkTop make b_compile
package Top(mkClkDivider, ClkDivider(..)) where

data State = IDLE | START | DATA (UInt (TLog 8)) | PARITY | STOP
  deriving (Bits, Eq, FShow)

type FCLK = 25_000_000
type BAUD = 9_600

interface (ClkDivider :: # -> *) hi =
  {
  reset :: Action
  ;isAdvancing :: Bool
  ;isHalfCycle :: Bool
  }

mkClkDivider :: Module (ClkDivider hi)
mkClkDivider = do
    counter <- mkReg(0 :: UInt (TLog hi))   
    let hi_value :: UInt (TLog hi) = (fromInteger $ valueOf hi)
    let half_hi_value :: UInt (TLog hi) = (fromInteger $ valueOf (TDiv hi 2))

    let val :: Real = (fromInteger $ valueOf hi)
    let msg = "Clock Div Period : " + (realToString val)
    -- messageM msg

    fileHandle <- openFile "compile.log" WriteMode 
    hPutStr fileHandle msg
    hClose fileHandle

    addRules $
      rules
        {-# ASSERT fire when enabled #-}
        {-# ASSERT no implicit conditions #-}
        "tick" : when True ==> action
          $display (counter)
          counter := if (counter == hi_value)
                    then 0
                    else counter + 1
    
    return $
      interface ClkDivider
        reset :: Action
        reset = do
          counter := 0

        isAdvancing :: Bool
        isAdvancing = (counter == hi_value)
        isHalfCycle = (counter == half_hi_value)

interface ITop = 
  ftdi_rxd    ::  Bit 1            {-# always_ready #-}
  led         ::  Bit 8            {-# always_ready #-}
  ftdi_txd    :: (Bit 1) -> Action {-# always_enabled, always_ready #-}

{-# properties mkTop={verilog} #-}
mkTop :: Module (ITop)
mkTop = do
  -- figure out why changing to wire below doesn't work
  ftdiRxIn :: Reg(Bit 1) <- mkReg(0)
  ledOutTemp :: Reg(Bit 8) <- mkReg(255)
  shiftReg :: Reg(Bit 8) <- mkReg(0)
  ftdiState <- mkReg(IDLE)

  clkDivider :: (ClkDivider (TDiv FCLK BAUD)) <- mkClkDivider

  addRules $
    rules

      {-# ASSERT fire when enabled #-}
      "exitIDLE" : when (ftdiState == IDLE), (ftdiRxIn == 0) ==>
        do
          clkDivider.reset
          ftdiState := START 

      {-# ASSERT fire when enabled #-}
      "exitSTART" : when (ftdiState == START), (clkDivider.isAdvancing) ==>
        do
          ftdiState := DATA(0)

      {-# ASSERT fire when enabled #-}
      "captureData" : 
        when 
          DATA(n) <- ftdiState,
          n >= 0,
          n <= 7, 
          let sampleTrigger = clkDivider.isHalfCycle
            in sampleTrigger
          ==>
            do
              ftdiState := 
                if n == 7
                  then PARITY
                  else DATA(n + 1)
              shiftReg := ftdiRxIn ++ shiftReg[7:1]

      {-# ASSERT fire when enabled #-}
      "exitPARITY" : when (ftdiState == PARITY), (clkDivider.isAdvancing) ==>
        do
          ftdiState := STOP

      {-# ASSERT fire when enabled #-}
      "exitSTOP" : when (ftdiState == STOP), (clkDivider.isAdvancing) ==>
        do
          ftdiState := IDLE

  return $
    interface ITop
    {led      = shiftReg
     ;ftdi_rxd = ftdiRxIn
     -- change below to do notation
     ;ftdi_txd bit = ftdiRxIn := bit
    }

mkSim :: Module Empty
mkSim = do
  -- count :: Reg(UInt 3) <- mkReg(0)
  count :: Reg(UInt 3) <- mkReg(0)
  addRules $
    rules
      "count" : when True ==> action
        count := unpack ((1'b1) ++ (pack count)[2:1])
        $display count
      "end sim" : when (count == 6) ==> action
        $finish

  return $
    interface Empty